module Memory_stage #(
    parameter D_WIDTH = 32,
    parameter A_WIDTH = 5
) (

);






endmodule
